--------------------------------------------------------------------------------
-- b8008_top_tb.vhdl
--------------------------------------------------------------------------------
-- Generic testbench for b8008_top - Complete system test
--
-- ROM-agnostic: Runs any program loaded via ROM_FILE generic
-- Outputs detailed register and state information for post-processing
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.b8008_types.all;

entity b8008_top_tb is
    generic (
        ROM_FILE : string := "test_programs/alu_test_as.mem"
    );
end entity b8008_top_tb;

architecture testbench of b8008_top_tb is

    -- Component declaration
    component b8008_top is
        generic (
            ROM_FILE : string := "test_programs/alu_test_as.mem"
        );
        port (
            clk_in      : in  std_logic;
            reset       : in  std_logic;
            interrupt   : in  std_logic;
            phi1_out    : out std_logic;
            phi2_out    : out std_logic;
            sync_out    : out std_logic;
            s0_out      : out std_logic;
            s1_out      : out std_logic;
            s2_out      : out std_logic;
            address_out : out std_logic_vector(13 downto 0);
            data_out    : out std_logic_vector(7 downto 0);
            ram_byte_0  : out std_logic_vector(7 downto 0);
            debug_reg_a         : out std_logic_vector(7 downto 0);
            debug_reg_b         : out std_logic_vector(7 downto 0);
            debug_reg_c         : out std_logic_vector(7 downto 0);
            debug_reg_d         : out std_logic_vector(7 downto 0);
            debug_reg_e         : out std_logic_vector(7 downto 0);
            debug_reg_h         : out std_logic_vector(7 downto 0);
            debug_reg_l         : out std_logic_vector(7 downto 0);
            debug_cycle         : out integer range 1 to 3;
            debug_pc            : out std_logic_vector(13 downto 0);
            debug_ir            : out std_logic_vector(7 downto 0);
            debug_needs_address : out std_logic;
            debug_int_pending   : out std_logic;
            debug_flag_carry    : out std_logic;
            debug_flag_zero     : out std_logic;
            debug_flag_sign     : out std_logic;
            debug_flag_parity   : out std_logic;
            debug_io_port_8     : out std_logic_vector(7 downto 0);
            debug_io_port_9     : out std_logic_vector(7 downto 0);
            debug_io_port_10    : out std_logic_vector(7 downto 0)
        );
    end component;

    -- Test signals
    signal clk_in      : std_logic := '0';
    signal reset       : std_logic := '1';
    signal interrupt   : std_logic := '0';
    signal phi1_out    : std_logic;
    signal phi2_out    : std_logic;
    signal sync_out    : std_logic;
    signal s0_out      : std_logic;
    signal s1_out      : std_logic;
    signal s2_out      : std_logic;
    signal address_out : std_logic_vector(13 downto 0);
    signal data_out    : std_logic_vector(7 downto 0);
    signal ram_byte_0  : std_logic_vector(7 downto 0);
    signal debug_reg_a         : std_logic_vector(7 downto 0);
    signal debug_reg_b         : std_logic_vector(7 downto 0);
    signal debug_reg_c         : std_logic_vector(7 downto 0);
    signal debug_reg_d         : std_logic_vector(7 downto 0);
    signal debug_reg_e         : std_logic_vector(7 downto 0);
    signal debug_reg_h         : std_logic_vector(7 downto 0);
    signal debug_reg_l         : std_logic_vector(7 downto 0);
    signal debug_cycle         : integer range 1 to 3;
    signal debug_pc            : std_logic_vector(13 downto 0);
    signal debug_ir            : std_logic_vector(7 downto 0);
    signal debug_needs_address : std_logic;
    signal debug_int_pending   : std_logic;
    signal debug_flag_carry    : std_logic;
    signal debug_flag_zero     : std_logic;
    signal debug_flag_sign     : std_logic;
    signal debug_flag_parity   : std_logic;
    signal debug_io_port_8     : std_logic_vector(7 downto 0);
    signal debug_io_port_9     : std_logic_vector(7 downto 0);
    signal debug_io_port_10    : std_logic_vector(7 downto 0);

    -- Clock generation
    constant CLK_PERIOD : time := 10 ns;  -- 100 MHz
    signal test_running : boolean := true;

    -- Test monitoring
    signal instruction_count : integer := 0;
    signal last_address : unsigned(13 downto 0) := (others => '0');
    signal stuck_counter : integer := 0;

begin

    -- ========================================================================
    -- DEVICE UNDER TEST
    -- ========================================================================

    dut : b8008_top
        generic map (
            ROM_FILE => ROM_FILE
        )
        port map (
            clk_in      => clk_in,
            reset       => reset,
            interrupt   => interrupt,
            phi1_out    => phi1_out,
            phi2_out    => phi2_out,
            sync_out    => sync_out,
            s0_out      => s0_out,
            s1_out      => s1_out,
            s2_out      => s2_out,
            address_out => address_out,
            data_out    => data_out,
            ram_byte_0  => ram_byte_0,
            debug_reg_a         => debug_reg_a,
            debug_reg_b         => debug_reg_b,
            debug_reg_c         => debug_reg_c,
            debug_reg_d         => debug_reg_d,
            debug_reg_e         => debug_reg_e,
            debug_reg_h         => debug_reg_h,
            debug_reg_l         => debug_reg_l,
            debug_cycle         => debug_cycle,
            debug_pc            => debug_pc,
            debug_ir            => debug_ir,
            debug_needs_address => debug_needs_address,
            debug_int_pending   => debug_int_pending,
            debug_flag_carry    => debug_flag_carry,
            debug_flag_zero     => debug_flag_zero,
            debug_flag_sign     => debug_flag_sign,
            debug_flag_parity   => debug_flag_parity,
            debug_io_port_8     => debug_io_port_8,
            debug_io_port_9     => debug_io_port_9,
            debug_io_port_10    => debug_io_port_10
        );

    -- ========================================================================
    -- CLOCK GENERATION
    -- ========================================================================

    clk_process : process
    begin
        while test_running loop
            clk_in <= '0';
            wait for CLK_PERIOD / 2;
            clk_in <= '1';
            wait for CLK_PERIOD / 2;
        end loop;
        wait;
    end process;

    -- ========================================================================
    -- STIMULUS AND MONITORING
    -- ========================================================================

    stimulus : process
    begin
        report "========================================";
        report "B8008 TOP-LEVEL SYSTEM TEST";
        report "Running search program from Intel 8008 User's Manual";
        report "========================================";

        -- Hold reset and interrupt low
        reset <= '1';
        interrupt <= '0';
        wait for 200 ns;

        -- Release reset
        reset <= '0';
        report "Reset released - CPU in stopped state";
        wait for 100 ns;

        -- Assert bootstrap interrupt to start CPU
        interrupt <= '1';
        wait for 1 ns;
        report "Bootstrap interrupt asserted";

        -- Wait for T1I state (S2='1', S1='1', S0='0'), then lower interrupt
        wait until (s2_out = '1' and s1_out = '1' and s0_out = '0');
        wait for 50 ns;  -- Wait a bit into T1I
        interrupt <= '0';
        report "T1I detected - interrupt lowered";
        wait for 100 ns;

        -- Let CPU run for a while and monitor execution
        report "Monitoring CPU execution...";

        -- Wait for CPU to execute the search program
        -- The program searches for '.' in "Hello, world. 8008!!"
        -- Expected: Program should find '.' at position 213 (0xD5) and halt

        -- Monitor for much longer to let program complete
        for i in 1 to 200000 loop
            wait for 100 ns;

            -- Report state periodically with debug info in clear format
            if i mod 100 = 0 then
                report "========================================";
                report "Cycle " & integer'image(i) & " @ " & time'image(now);
                report "  PC = 0x" & to_hstring(unsigned(debug_pc)) &
                       " | IR = 0x" & to_hstring(unsigned(debug_ir)) &
                       " | MCycle = " & integer'image(debug_cycle);
                report "CPU Registers (scratchpad):";
                report "  Reg.A = 0x" & to_hstring(unsigned(debug_reg_a)) &
                       " | Reg.B = 0x" & to_hstring(unsigned(debug_reg_b)) &
                       " | Reg.C = 0x" & to_hstring(unsigned(debug_reg_c));
                report "  Reg.D = 0x" & to_hstring(unsigned(debug_reg_d)) &
                       " | Reg.E = 0x" & to_hstring(unsigned(debug_reg_e));
                report "  Reg.H = 0x" & to_hstring(unsigned(debug_reg_h)) &
                       " | Reg.L = 0x" & to_hstring(unsigned(debug_reg_l)) &
                       "  (H:L ptr = " & integer'image(to_integer(unsigned(debug_reg_h & debug_reg_l))) & ")";
                report "Flags: C=" & std_logic'image(debug_flag_carry) &
                       " Z=" & std_logic'image(debug_flag_zero) &
                       " S=" & std_logic'image(debug_flag_sign) &
                       " P=" & std_logic'image(debug_flag_parity);
                report "External Bus:";
                report "  Addr = 0x" & to_hstring(unsigned(address_out)) &
                       " | Data = 0x" & to_hstring(unsigned(data_out)) &
                       " | State = " & std_logic'image(s2_out) &
                       std_logic'image(s1_out) & std_logic'image(s0_out);
            end if;

            -- Check if address changed (new instruction fetch)
            if unsigned(address_out) /= last_address then
                last_address <= unsigned(address_out);

                -- Report all addresses for first 50us to debug
                if now < 50 us then
                    report "  @" & time'image(now) & " Addr=0x" & to_hstring(unsigned(address_out)) &
                           " Data=0x" & to_hstring(unsigned(data_out)) &
                           " State=" & std_logic'image(s2_out) & std_logic'image(s1_out) & std_logic'image(s0_out);
                end if;

                -- Report key addresses
                if address_out = x"0000" then
                    report "  ** Fetching from 0x0000 (Reset vector)";
                elsif address_out = x"0100" then
                    report "  ** Reached MAIN at 0x0100";
                elsif address_out = x"003C" then
                    report "  ** Calling INCR subroutine at 0x003C";
                elsif unsigned(address_out) >= 200 and unsigned(address_out) <= 220 then
                    report "  ** Reading string data at 0x" & to_hstring(unsigned(address_out)) &
                           " = '" & character'val(to_integer(unsigned(data_out))) & "'";
                end if;
            end if;

            -- Removed halt detection logic - was misleading during debugging
        end loop;

        wait for 1 us;

        report "========================================";
        report "SIMULATION COMPLETE";
        report "========================================";
        report "Simulation time: 20ms";
        report " ";
        report "Use external verification scripts to validate results.";
        report "Output above contains cycle-by-cycle register state.";
        report "========================================";

        -- End simulation
        test_running <= false;
        wait;
    end process;

end architecture testbench;
