--------------------------------------------------------------------------------
-- program_counter.vhdl
--------------------------------------------------------------------------------
-- Simple, explicit program counter for Intel 8008
--
-- This module does ONE thing: manages the 14-bit program counter
-- - Increments when increment control is high (level-triggered latch)
-- - Loads when load control is high (level-triggered latch)
-- - Holds when hold control is high or all controls low
-- - NO clock signal - uses level-triggered latches (1972 design)
-- - NO conditional logic, NO knowledge of instructions or interrupts
--
-- Note: Control signals are pulses/strobes generated by timing/control logic
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.b8008_types.all;

entity program_counter is
    port (
        -- Control signals (explicit, one-hot pulses/strobes)
        control   : in  pc_control_t;

        -- Data input for load operation
        data_in   : in  address_t;

        -- Current PC value (always available)
        pc_out    : out address_t
    );
end entity program_counter;

architecture rtl of program_counter is
    signal pc : address_t := (others => '0');
begin

    -- Output current PC
    pc_out <= pc;

    -- Latch behavior: respond to rising edge of control strobes
    -- In real 1972 hardware, these would be level-triggered latches
    -- In VHDL simulation, we model the strobe edge to avoid delta cycles
    process(control.increment, control.load)
    begin
        -- Increment on rising edge of increment strobe
        if rising_edge(control.increment) then
            pc <= pc + 1;

        -- Load on rising edge of load strobe
        elsif rising_edge(control.load) then
            pc <= data_in;
        end if;

        -- Hold is implicit - no edge means no change
    end process;

end architecture rtl;
