-------------------------------------------------------------------------------
-- Intel 8008 v8008 INP (Input from Port) Instruction Test
-------------------------------------------------------------------------------
-- Tests INP instruction (opcode 0x41-0x4F, pattern: 01 00M MM1):
-- - Reads data from one of 8 input ports (MMM = 0-7) into accumulator
-- - Two-cycle instruction (fetch + I/O read)
-- - Cycle 0: Standard instruction fetch
-- - Cycle 1: 5-state I/O cycle (T1-T5) with PCC cycle type
-- - Verifies accumulator receives I/O data
-- - Verifies flag output at T4
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use STD.TEXTIO.ALL;

entity v8008_inp_tb is
end v8008_inp_tb;

architecture behavior of v8008_inp_tb is

    -- Component declaration for v8008 CPU
    component v8008
        port (
            -- Two-phase clock inputs
            phi1 : in std_logic;
            phi2 : in std_logic;

            -- Data bus
            data_bus_in     : in  std_logic_vector(7 downto 0);
            data_bus_out    : out std_logic_vector(7 downto 0);
            data_bus_enable : out std_logic;

            -- State outputs
            S0 : out std_logic;
            S1 : out std_logic;
            S2 : out std_logic;

            -- SYNC output
            SYNC : out std_logic;

            -- READY input
            READY : in std_logic;

            -- Interrupt request
            INT : in std_logic;

            -- Debug outputs
            debug_reg_A : out std_logic_vector(7 downto 0);
            debug_reg_B : out std_logic_vector(7 downto 0);
            debug_reg_C : out std_logic_vector(7 downto 0);
            debug_reg_D : out std_logic_vector(7 downto 0);
            debug_reg_E : out std_logic_vector(7 downto 0);
            debug_reg_H : out std_logic_vector(7 downto 0);
            debug_reg_L : out std_logic_vector(7 downto 0);
            debug_pc : out std_logic_vector(13 downto 0);
            debug_flags : out std_logic_vector(3 downto 0);
            debug_instruction : out std_logic_vector(7 downto 0);
            debug_stack_pointer : out std_logic_vector(2 downto 0);
            debug_hl_address : out std_logic_vector(13 downto 0)
        );
    end component;

    -- Clock and control signals
    signal phi1        : std_logic := '0';
    signal phi2        : std_logic := '0';
    signal INT         : std_logic := '0';
    signal READY       : std_logic := '1';

    -- CPU interface
    signal data_bus_in : std_logic_vector(7 downto 0) := (others => '0');
    signal data_bus_out: std_logic_vector(7 downto 0);
    signal data_bus_enable : std_logic;
    signal S0          : std_logic;
    signal S1          : std_logic;
    signal S2          : std_logic;
    signal SYNC        : std_logic;

    -- Debug signals
    signal debug_reg_A : std_logic_vector(7 downto 0);
    signal debug_reg_B : std_logic_vector(7 downto 0);
    signal debug_reg_C : std_logic_vector(7 downto 0);
    signal debug_reg_D : std_logic_vector(7 downto 0);
    signal debug_reg_E : std_logic_vector(7 downto 0);
    signal debug_reg_H : std_logic_vector(7 downto 0);
    signal debug_reg_L : std_logic_vector(7 downto 0);
    signal debug_pc    : std_logic_vector(13 downto 0);
    signal debug_flags : std_logic_vector(3 downto 0);
    signal debug_instruction : std_logic_vector(7 downto 0);
    signal debug_stack_pointer : std_logic_vector(2 downto 0);
    signal debug_hl_address : std_logic_vector(13 downto 0);

    -- Test control
    signal done        : boolean := false;
    signal test_phase  : string(1 to 20) := (others => ' ');
    signal test_num    : integer := 0;

    -- Constants
    constant PHI1_PERIOD : time := 1100 ns;
    constant PHI2_PERIOD : time := 1100 ns;
    constant OVERLAP_TIME : time := 100 ns;

    -- Test cases for INP instruction
    type test_case_t is record
        port_num : integer range 0 to 7;        -- Port number (MMM bits)
        opcode   : std_logic_vector(7 downto 0);  -- INP opcode
        io_data  : std_logic_vector(7 downto 0);  -- Data to provide from I/O port
        description : string(1 to 30);
    end record;

    type test_cases_array_t is array (0 to 7) of test_case_t;
    constant test_cases : test_cases_array_t := (
        -- Test all 8 input ports with different data patterns
        (port_num => 0, opcode => x"41", io_data => x"AA", description => "INP Port 0, data 0xAA         "),
        (port_num => 1, opcode => x"43", io_data => x"55", description => "INP Port 1, data 0x55         "),
        (port_num => 2, opcode => x"45", io_data => x"FF", description => "INP Port 2, data 0xFF         "),
        (port_num => 3, opcode => x"47", io_data => x"00", description => "INP Port 3, data 0x00         "),
        (port_num => 4, opcode => x"49", io_data => x"42", description => "INP Port 4, data 0x42         "),
        (port_num => 5, opcode => x"4B", io_data => x"CC", description => "INP Port 5, data 0xCC         "),
        (port_num => 6, opcode => x"4D", io_data => x"33", description => "INP Port 6, data 0x33         "),
        (port_num => 7, opcode => x"4F", io_data => x"F0", description => "INP Port 7, data 0xF0         ")
    );

    -- I/O simulation
    signal current_port : integer range 0 to 7 := 0;
    signal io_port_data : std_logic_vector(7 downto 0) := x"00";

    -- Cycle tracking for I/O detection
    signal cpu_cycle : integer range 0 to 2 := 0;
    signal prev_state : std_logic_vector(2 downto 0) := "011";  -- Start at STOPPED

begin

    -- Instantiate v8008 CPU
    UUT: v8008
        port map (
            phi1 => phi1,
            phi2 => phi2,
            data_bus_in => data_bus_in,
            data_bus_out => data_bus_out,
            data_bus_enable => data_bus_enable,
            S0 => S0,
            S1 => S1,
            S2 => S2,
            SYNC => SYNC,
            READY => READY,
            INT => INT,
            debug_reg_A => debug_reg_A,
            debug_reg_B => debug_reg_B,
            debug_reg_C => debug_reg_C,
            debug_reg_D => debug_reg_D,
            debug_reg_E => debug_reg_E,
            debug_reg_H => debug_reg_H,
            debug_reg_L => debug_reg_L,
            debug_pc => debug_pc,
            debug_flags => debug_flags,
            debug_instruction => debug_instruction,
            debug_stack_pointer => debug_stack_pointer,
            debug_hl_address => debug_hl_address
        );

    -- Cycle tracking process
    CYCLE_TRACK: process
        variable state_vec : std_logic_vector(2 downto 0);
        variable instr_complete : boolean;
    begin
        wait on S0, S1, S2, debug_instruction;
        state_vec := S2 & S1 & S0;

        -- Determine if instruction is complete based on debug_instruction
        -- HLT doesn't transition to another instruction, but INP does
        instr_complete := ((debug_instruction(7 downto 6) = "01" and
                           debug_instruction(5 downto 4) = "00" and
                           debug_instruction(0) = '1') or  -- INP instruction
                          (debug_instruction /= x"00" and debug_instruction /= x"FF"));  -- Not HLT

        -- Track cycle transitions
        if state_vec = "011" then  -- STOPPED - reset cycle
            cpu_cycle <= 0;
        elsif state_vec = "110" then  -- T1I - always cycle 0 (interrupt ack)
            cpu_cycle <= 0;
        elsif (prev_state = "001" or prev_state = "101") and state_vec = "010" then  -- T3/T5 -> T1
            -- Check if this is a new instruction (cycle increment) or new cycle
            -- For multi-cycle instructions, increment cycle
            -- For instruction completion, reset to 0
            if cpu_cycle = 1 and instr_complete then
                cpu_cycle <= 0;  -- Instruction complete, start next instruction at cycle 0
            elsif cpu_cycle < 2 then
                cpu_cycle <= cpu_cycle + 1;  -- Multi-cycle instruction, increment
            end if;
        end if;

        prev_state <= state_vec;
    end process CYCLE_TRACK;

    -- Memory and I/O simulation process
    MEM_IO_PROC: process
        variable state_vec : std_logic_vector(2 downto 0);
        variable decoded_port : integer range 0 to 7;
        variable is_inp_instruction : boolean;
    begin
        wait on S0, S1, S2, data_bus_out, data_bus_enable, cpu_cycle, debug_instruction;

        state_vec := S2 & S1 & S0;

        -- Check if current instruction is INP
        is_inp_instruction := (debug_instruction(7 downto 6) = "01" and
                              debug_instruction(5 downto 4) = "00" and
                              debug_instruction(0) = '1');

        -- Handle operations based on state
        case state_vec is
            when "001" =>  -- T3: Data transfer state
                -- Check if CPU is driving the bus or expecting input
                if data_bus_enable = '0' then
                    -- CPU is reading - determine what to provide
                    -- Check if we're in cycle 1 of an INP instruction (I/O read)
                    if cpu_cycle = 1 and is_inp_instruction then
                        -- I/O read - decode port from instruction and provide corresponding data
                        decoded_port := to_integer(unsigned(debug_instruction(3 downto 1)));
                        data_bus_in <= test_cases(decoded_port).io_data;
                        report "I/O: Providing data 0x" & to_hstring(test_cases(decoded_port).io_data) &
                               " from port " & integer'image(decoded_port) &
                               " (cycle=" & integer'image(cpu_cycle) & ")";
                    elsif to_integer(unsigned(debug_pc)) < 100 then
                        -- Program area - provide instructions
                        -- Sequential INP instructions (no HLT between them)
                        case to_integer(unsigned(debug_pc)) is
                            when 0  => data_bus_in <= test_cases(0).opcode;  -- INP port 0
                            when 1  => data_bus_in <= test_cases(1).opcode;  -- INP port 1
                            when 2  => data_bus_in <= test_cases(2).opcode;  -- INP port 2
                            when 3  => data_bus_in <= test_cases(3).opcode;  -- INP port 3
                            when 4  => data_bus_in <= test_cases(4).opcode;  -- INP port 4
                            when 5  => data_bus_in <= test_cases(5).opcode;  -- INP port 5
                            when 6  => data_bus_in <= test_cases(6).opcode;  -- INP port 6
                            when 7  => data_bus_in <= test_cases(7).opcode;  -- INP port 7
                            when 8  => data_bus_in <= x"FF";  -- HLT at end

                            when others => data_bus_in <= x"FF";  -- HLT
                        end case;
                    else
                        -- Default
                        data_bus_in <= x"00";
                    end if;
                end if;

            when "111" =>  -- T4: Flag output for I/O
                -- CPU should be driving flags during INP
                if data_bus_enable = '1' then
                    report "T4: Flags output detected: 0x" & to_hstring(data_bus_out);
                end if;

            when others =>
                -- Other states - provide default
                null;
        end case;
    end process MEM_IO_PROC;

    -- Clock generation
    CLOCK_PROC: process
    begin
        while not done loop
            -- phi1 high phase
            phi1 <= '1';
            wait for PHI1_PERIOD - OVERLAP_TIME;

            -- phi2 rises while phi1 still high (overlap)
            phi2 <= '1';
            wait for OVERLAP_TIME;

            -- phi1 falls, phi2 stays high
            phi1 <= '0';
            wait for PHI2_PERIOD - OVERLAP_TIME;

            -- phi2 falls
            phi2 <= '0';
            wait for OVERLAP_TIME;
        end loop;
        wait;
    end process CLOCK_PROC;

    -- Main test process
    TEST_PROC: process
        variable state_vec : std_logic_vector(2 downto 0);
        variable initial_pc : std_logic_vector(13 downto 0);
        variable initial_acc : std_logic_vector(7 downto 0);
    begin
        report "========================================";
        report "Intel 8008 INP Instruction Test";
        report "Testing Input from Port (0x41-0x4F)";
        report "========================================";

        -- Initialize CPU (trigger interrupt to start from known state)
        test_phase <= "INIT                ";
        wait for 500 ns;

        -- CPU starts in STOPPED state
        state_vec := S2 & S1 & S0;
        assert state_vec = "011"
            report "ERROR: CPU not starting in STOPPED state"
            severity error;

        -- Trigger interrupt once to start CPU
        report "";
        report "Starting CPU execution...";
        wait until rising_edge(phi1);
        INT <= '1';
        wait for 3000 ns;
        INT <= '0';

        -- Test each INP instruction for all 8 ports
        -- They execute sequentially without interrupts
        for i in 0 to 7 loop
            test_num <= i;

            case i is
                when 0 => test_phase <= "TEST 0              ";
                when 1 => test_phase <= "TEST 1              ";
                when 2 => test_phase <= "TEST 2              ";
                when 3 => test_phase <= "TEST 3              ";
                when 4 => test_phase <= "TEST 4              ";
                when 5 => test_phase <= "TEST 5              ";
                when 6 => test_phase <= "TEST 6              ";
                when 7 => test_phase <= "TEST 7              ";
                when others => test_phase <= "TEST ?              ";
            end case;

            report "";
            report "Test " & integer'image(i + 1) & ": " & test_cases(i).description;
            report "  Port = " & integer'image(test_cases(i).port_num);
            report "  Opcode = 0x" & to_hstring(test_cases(i).opcode);
            report "  I/O Data = 0x" & to_hstring(test_cases(i).io_data);
            report "--------------------------------------";

            -- Wait for INP instruction to complete
            -- Each INP: Cycle 0 (~7us) + Cycle 1 (~11us) = ~18us
            wait for 20000 ns;

            -- Verify accumulator received I/O data
            assert debug_reg_A = test_cases(i).io_data
                report "ERROR: Accumulator did not receive I/O data. Expected 0x" &
                       to_hstring(test_cases(i).io_data) &
                       ", got 0x" & to_hstring(debug_reg_A)
                severity error;

            report "Accumulator after INP: 0x" & to_hstring(debug_reg_A) & " (correct)";
            report "PASS: INP test " & integer'image(i + 1) & " successful";
        end loop;

        -- Wait for HLT at the end
        wait for 10000 ns;
        state_vec := S2 & S1 & S0;
        assert state_vec = "011"
            report "WARNING: CPU not in STOPPED state after final HLT"
            severity warning;

        ------------------------------
        -- Test complete
        ------------------------------
        test_phase <= "DONE                ";
        report "";
        report "========================================";
        report "INP Test Summary:";
        report "  - All 8 input ports tested: PASS";
        report "  - Opcode fetch and PC increment: PASS";
        report "  - I/O data transfer to accumulator: PASS";
        report "  - 2-cycle I/O operation timing: PASS";
        report "========================================";

        done <= true;
        wait;
    end process TEST_PROC;

end behavior;
